// This is the parameter definition for the VP unit
//
`define VP_ENABLED
`define P_CONF_WIDTH 8
`define P_STORAGE_SIZE 2048