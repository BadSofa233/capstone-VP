03CE0E3300100E13
03CE0E3303CE0E33
FE0008E303CE0E33
0000000000000013
