006E0E1300000E13
003E7E13FFFE0E13
00000013FE000AE3
0000000000000000
